// Copyright (C) 2022  The Symbiflow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC

module top (
    input  wire clk,

    input  wire rx,
    output wire tx,

    input  wire [15:0] sw,
    output wire [15:0] led
);
    RAM64M8 #(
        // FIXME: python-fpga_interchange seems to be unable to parse any literal wider than 64-bit
        //.INIT_A(128'b10101010101010101010101010101010101010101010101010101010101010100000000111111111111111011111100111110001111000011100000110000001),
        //.INIT_B(128'b11001100110011001100110011001100110011001100110011001100110011000000001111111111111110111111001111100011110000111000001100000010),
        //.INIT_C(128'b11110000111100001111000011110000111100001111000011110000111100000000011111111111111101111110011111000111100001110000011000000100),
        //.INIT_D(128'b11111111000000001111111100000000111111110000000011111111000000000000111111111111111011111100111110001111000011100000110000001000),
        //.INIT_E(128'b11111111111111110000000000000000111111111111111100000000000000000001111111111111110111111001111100011110000111000001100000010000),
        //.INIT_F(128'b11111111111111111111111111111111000000000000000000000000000000000011111111111111101111110011111000111100001110000011000000100000),
        //.INIT_G(128'b10110011100011110000111110000011111100000011111110000000111111110111111111111111011111100111110001111000011100000110000001000000),
        //.INIT_H(128'b01001100011100001111000001111100000011111100000001111111000000001111111111111110111111001111100011110000111000001100000010000000)
        .INIT_A(128'b0000000111111111111111011111100111110001111000011100000110000001),
        .INIT_B(128'b0000001111111111111110111111001111100011110000111000001100000010),
        .INIT_C(128'b0000011111111111111101111110011111000111100001110000011000000100),
        .INIT_D(128'b0000111111111111111011111100111110001111000011100000110000001000),
        .INIT_E(128'b0001111111111111110111111001111100011110000111000001100000010000),
        .INIT_F(128'b0011111111111111101111110011111000111100001110000011000000100000),
        .INIT_G(128'b0111111111111111011111100111110001111000011100000110000001000000),
        .INIT_H(128'b1111111111111110111111001111100011110000111000001100000010000000)
    ) ram0 (
        .WCLK   (clk),
        .ADDRA  (sw[5:0]),
        .ADDRB  (sw[5:0]),
        .ADDRC  (sw[5:0]),
        .ADDRD  (sw[5:0]),
        .ADDRE  (sw[5:0]),
        .ADDRF  (sw[5:0]),
        .ADDRG  (sw[5:0]),
        .ADDRH  (sw[5:0]),
        .DIA    (sw[12]),
        .DIB    (sw[13]),
        .DIC    (sw[14]),
        .DID    (sw[14]),
        .DID    (sw[14]),
        .DID    (sw[14]),
        .DID    (sw[14]),
        .DID    (sw[14]),
        .DOA    (led[0]),
        .DOB    (led[1]),
        .DOC    (led[2]),
        .DOD    (led[3]),
        .WE     (sw[15])
    );

    assign led[15:8] = sw[15:8];
    assign tx = rx;

endmodule
