// Copyright (C) 2021  The Symbiflow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC

// Inverter support is still a TODO
module INV(input A, output Z);
	LUT4 #(.INIT("0x5555")) _TECHMAP_REPLACE_ (.A(A), .B(1'b1), .C(1'b1), .D(1'b1), .Z(Z));
endmodule

module PDPSC16K (...);
	parameter DATA_WIDTH_W = "X36";
	parameter DATA_WIDTH_R = "X36";
	parameter OUTREG = "BYPASSED";
	parameter RESETMODE = "SYNC";
	parameter GSR = "ENABLED";
	parameter ECC = "DISABLED";
	parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
	parameter CSDECODE_W = "000";
	parameter CSDECODE_R = "000";
	parameter ASYNC_RST_RELEASE = "SYNC";
	parameter INIT_DATA = "STATIC";
	input [35:0] DI;
	input [13:0] ADW;
	input [13:0] ADR;
	input CLK;
	input CER;
	input CEW;
	input [2:0] CSW;
	input [2:0] CSR;
	input RST;
	output [35:0] DO;
	output ONEBITERR;
	output TWOBITERR;

	// TODO: this should really be a macro or otherwise dealt with more automatically
	PDPSC16K_MODE #(
		.DATA_WIDTH_W(DATA_WIDTH_W),
		.DATA_WIDTH_R(DATA_WIDTH_R),
		.OUTREG(OUTREG),
		.GSR(GSR),
		.ECC(ECC),
		.CSDECODE_W(CSDECODE_W),
		.CSDECODE_R(CSDECODE_R),
		.ASYNC_RST_RELEASE(ASYNC_RST_RELEASE),
		.INITVAL_00(INITVAL_00),
		.INITVAL_01(INITVAL_01),
		.INITVAL_02(INITVAL_02),
		.INITVAL_03(INITVAL_03),
		.INITVAL_04(INITVAL_04),
		.INITVAL_05(INITVAL_05),
		.INITVAL_06(INITVAL_06),
		.INITVAL_07(INITVAL_07),
		.INITVAL_08(INITVAL_08),
		.INITVAL_09(INITVAL_09),
		.INITVAL_0A(INITVAL_0A),
		.INITVAL_0B(INITVAL_0B),
		.INITVAL_0C(INITVAL_0C),
		.INITVAL_0D(INITVAL_0D),
		.INITVAL_0E(INITVAL_0E),
		.INITVAL_0F(INITVAL_0F),
		.INITVAL_10(INITVAL_10),
		.INITVAL_11(INITVAL_11),
		.INITVAL_12(INITVAL_12),
		.INITVAL_13(INITVAL_13),
		.INITVAL_14(INITVAL_14),
		.INITVAL_15(INITVAL_15),
		.INITVAL_16(INITVAL_16),
		.INITVAL_17(INITVAL_17),
		.INITVAL_18(INITVAL_18),
		.INITVAL_19(INITVAL_19),
		.INITVAL_1A(INITVAL_1A),
		.INITVAL_1B(INITVAL_1B),
		.INITVAL_1C(INITVAL_1C),
		.INITVAL_1D(INITVAL_1D),
		.INITVAL_1E(INITVAL_1E),
		.INITVAL_1F(INITVAL_1F),
		.INITVAL_20(INITVAL_20),
		.INITVAL_21(INITVAL_21),
		.INITVAL_22(INITVAL_22),
		.INITVAL_23(INITVAL_23),
		.INITVAL_24(INITVAL_24),
		.INITVAL_25(INITVAL_25),
		.INITVAL_26(INITVAL_26),
		.INITVAL_27(INITVAL_27),
		.INITVAL_28(INITVAL_28),
		.INITVAL_29(INITVAL_29),
		.INITVAL_2A(INITVAL_2A),
		.INITVAL_2B(INITVAL_2B),
		.INITVAL_2C(INITVAL_2C),
		.INITVAL_2D(INITVAL_2D),
		.INITVAL_2E(INITVAL_2E),
		.INITVAL_2F(INITVAL_2F),
		.INITVAL_30(INITVAL_30),
		.INITVAL_31(INITVAL_31),
		.INITVAL_32(INITVAL_32),
		.INITVAL_33(INITVAL_33),
		.INITVAL_34(INITVAL_34),
		.INITVAL_35(INITVAL_35),
		.INITVAL_36(INITVAL_36),
		.INITVAL_37(INITVAL_37),
		.INITVAL_38(INITVAL_38),
		.INITVAL_39(INITVAL_39),
		.INITVAL_3A(INITVAL_3A),
		.INITVAL_3B(INITVAL_3B),
		.INITVAL_3C(INITVAL_3C),
		.INITVAL_3D(INITVAL_3D),
		.INITVAL_3E(INITVAL_3E),
		.INITVAL_3F(INITVAL_3F),
		.INIT_DATA(INIT_DATA)
	) _TECHMAP_REPLACE_ (
		.CLK(CLK), .CER(CER), .CEW(CEW), .RST(RST),
		.CSW0(CSW[0]), .CSW1(CSW[1]), .CSW2(CSW[2]),
		.CSR0(CSR[0]), .CSR1(CSR[1]), .CSR2(CSR[2]),
		.DI0(DI[0]), .DI1(DI[1]), .DI2(DI[2]), .DI3(DI[3]), .DI4(DI[4]), .DI5(DI[5]), .DI6(DI[6]), .DI7(DI[7]), .DI8(DI[8]), .DI9(DI[9]), .DI10(DI[10]), .DI11(DI[11]), .DI12(DI[12]), .DI13(DI[13]), .DI14(DI[14]), .DI15(DI[15]), .DI16(DI[16]), .DI17(DI[17]), .DI18(DI[18]), .DI19(DI[19]), .DI20(DI[20]), .DI21(DI[21]), .DI22(DI[22]), .DI23(DI[23]), .DI24(DI[24]), .DI25(DI[25]), .DI26(DI[26]), .DI27(DI[27]), .DI28(DI[28]), .DI29(DI[29]), .DI30(DI[30]), .DI31(DI[31]), .DI32(DI[32]), .DI33(DI[33]), .DI34(DI[34]), .DI35(DI[35]),
		.ADW0(ADW[0]), .ADW1(ADW[1]), .ADW2(ADW[2]), .ADW3(ADW[3]), .ADW4(ADW[4]), .ADW5(ADW[5]), .ADW6(ADW[6]), .ADW7(ADW[7]), .ADW8(ADW[8]), .ADW9(ADW[9]), .ADW10(ADW[10]), .ADW11(ADW[11]), .ADW12(ADW[12]), .ADW13(ADW[13]),
		.ADR0(ADR[0]), .ADR1(ADR[1]), .ADR2(ADR[2]), .ADR3(ADR[3]), .ADR4(ADR[4]), .ADR5(ADR[5]), .ADR6(ADR[6]), .ADR7(ADR[7]), .ADR8(ADR[8]), .ADR9(ADR[9]), .ADR10(ADR[10]), .ADR11(ADR[11]), .ADR12(ADR[12]), .ADR13(ADR[13]),
		.DO0(DO[0]), .DO1(DO[1]), .DO2(DO[2]), .DO3(DO[3]), .DO4(DO[4]), .DO5(DO[5]), .DO6(DO[6]), .DO7(DO[7]), .DO8(DO[8]), .DO9(DO[9]), .DO10(DO[10]), .DO11(DO[11]), .DO12(DO[12]), .DO13(DO[13]), .DO14(DO[14]), .DO15(DO[15]), .DO16(DO[16]), .DO17(DO[17]), .DO18(DO[18]), .DO19(DO[19]), .DO20(DO[20]), .DO21(DO[21]), .DO22(DO[22]), .DO23(DO[23]), .DO24(DO[24]), .DO25(DO[25]), .DO26(DO[26]), .DO27(DO[27]), .DO28(DO[28]), .DO29(DO[29]), .DO30(DO[30]), .DO31(DO[31]), .DO32(DO[32]), .DO33(DO[33]), .DO34(DO[34]), .DO35(DO[35]),
		.ONEBITERR(ONEBITERR), .TWOBITERR(TWOBITERR),
	);

endmodule
