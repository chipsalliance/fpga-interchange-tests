// Copyright (C) 2022  The Symbiflow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC

module top (
    input  wire clk,

    input  wire rx,
    output wire tx,

    input  wire [15:0] sw,
    output wire [15:0] led
);
    RAM32M16 #(
        // FIXME: python-fpga_interchange seems to be unable to parse any literal wider than 64-bit
        //.INIT_A(128'b00_00_00_00_00_00_00_00_00_00_00_00_00_00_10_11_11_11_01_00_00_00_00_00_00_00_00_00_00_00_10_11_11_01_00_00_00_00_00_00_00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01),
        //.INIT_B(128'b00_00_00_00_00_00_00_00_00_00_00_00_10_11_11_11_01_00_00_00_00_00_00_00_00_00_00_00_10_11_11_01_00_00_00_00_00_00_00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00),
        //.INIT_C(128'b00_00_00_00_00_00_00_00_00_00_10_11_11_11_01_00_00_00_00_00_00_00_00_00_00_00_10_11_11_01_00_00_00_00_00_00_00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00_00_00),
        //.INIT_D(128'b00_00_00_00_00_00_00_00_10_11_11_11_01_00_00_00_00_00_00_00_00_00_00_00_10_11_11_01_00_00_00_00_00_00_00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00_00_00_00_00),
        //.INIT_E(128'b00_00_00_00_00_00_10_11_11_11_01_00_00_00_00_00_00_00_00_00_00_00_10_11_11_01_00_00_00_00_00_00_00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00_00_00_00_00_00_00),
        //.INIT_F(128'b00_00_00_00_10_11_11_11_01_00_00_00_00_00_00_00_00_00_00_00_10_11_11_01_00_00_00_00_00_00_00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00_00_00_00_00_00_00_00_00),
        //.INIT_G(128'b00_00_10_11_11_11_01_00_00_00_00_00_00_00_00_00_00_00_10_11_11_01_00_00_00_00_00_00_00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00_00_00_00_00_00_00_00_00_00_00),
        //.INIT_H(128'b10_11_11_11_01_00_00_00_00_00_00_00_00_00_00_00_10_11_11_01_00_00_00_00_00_00_00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00_00_00_00_00_00_00_00_00_00_00_00_00)
        .INIT_A(128'b00_00_00_00_00_00_00_00_00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01),
        .INIT_B(128'b00_00_00_00_00_00_00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00),
        .INIT_C(128'b00_00_00_00_00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00_00_00),
        .INIT_D(128'b00_00_00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00_00_00_00_00),
        .INIT_E(128'b00_00_00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00_00_00_00_00_00_00),
        .INIT_F(128'b00_00_00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00_00_00_00_00_00_00_00_00),
        .INIT_G(128'b00_00_10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00_00_00_00_00_00_00_00_00_00_00),
        .INIT_H(128'b10_11_01_00_00_00_00_00_00_00_00_00_00_00_00_00_10_01_00_00_00_00_00_00_00_00_00_00_00_00_00_00)
    ) ram0 (
        .WCLK    (clk),
        .ADDRA   (sw[4:0]),
        .ADDRB   (sw[4:0]),
        .ADDRC   (sw[4:0]),
        .ADDRD   (sw[4:0]),
        .ADDRE   (sw[4:0]),
        .ADDRF   (sw[4:0]),
        .ADDRG   (sw[4:0]),
        .ADDRH   (sw[4:0]),
        .DIA     (sw[9:8]),
        .DIB     (sw[11:10]),
        .DIC     (sw[13:12]),
        .DID     (sw[15:14]),
        .DIE     (sw[11:10]),
        .DIF     (sw[11:10]),
        .DIG     (sw[13:12]),
        .DIH     (sw[15:14]),
        .DOA     (led[1:0]),
        .DOB     (led[3:2]),
        .DOC     (led[5:4]),
        .DOD     (led[7:6]),
        .DOE     (led[9:8]),
        .DOF     (led[11:10]),
        .DOG     (led[13:12]),
        .DOH     (led[15:14]),
        .WE      (sw[15])
    );

    assign tx = rx;

endmodule
